// Code your design here
module sync_fifo #(parameter width=8,parameter depth=8)(

input clk,
input rst,
input wr_en,
input rd_en,
input [width-1:0]data_in,
output reg [width-1:0] data_out,
output full,
output empty);
  
  //reg tflag;
              
reg [$clog2(depth):0]wr_ptr;
reg [$clog2(depth):0]rd_ptr;
  integer i;
  
  reg[width-1:0] fifo [depth-1:0];
  
  always@(posedge clk or negedge rst)
    begin 
      if(!rst)
        begin
          wr_ptr<=0;
          rd_ptr<=0;
//           empty<=1;
//           full<=0;
          
          for(i=0;i<depth;i=i+1)
            begin
              fifo[i]<=0;
            end
          
        end
      
      else 
        begin
        if(wr_en && !full)
        begin
          fifo[wr_ptr[$clog2(depth)-1:0]]<=data_in;
          wr_ptr<=wr_ptr+1;
          
         /* if(wr_ptr==fifo_depth-1)
            tflag<=1;*/
          
        end
      
       if(rd_en && !empty)
        begin
          data_out<=fifo[rd_ptr[$clog2(depth)-1:0]];
          rd_ptr<=rd_ptr+1;
      
        end
      
     
      
    end
    end
      //assign  empty= !rst ? 1'b1 :((wr_ptr==rd_ptr) && (tflag!=1));
      assign  empty= (wr_ptr==rd_ptr);
      assign full={~wr_ptr[$clog2(depth)],wr_ptr[$clog2(depth)-1:0]}==rd_ptr;
endmodule
